/**
* Costa Rica Institute of Technology
* @author Kendall González
* Computer Architecture
* ASIP
*/


// This file will be included in the other system verilog components
// will allow the change of the processor parameters easily

`define ALUSize 32 // size of the operands in bits that can handle the ALU
`define RegisterSize 32 // register's size in bits
`define AmountOfRegisters 16 // quantity of registers in the processor
`define ImageWidth 320 // Canvas size
`define ImageHeigth 240 // Canvas size
